module CORE(
  input CLK, RST
);

wire ALU, BRA, COND_BRA, BRZ, BRN, BRC, BRO, LOAD, STORE, COPY, PUSH, POP, MOV, SEL_FLAG, SEL_ACC, SEL_X, SEL_Y, SEL_PC;
wire [15:0] PC_VAL;
wire signed [15:0] ACC_VAL;
wire signed [15:0] X_VAL;
wire signed [15:0] Y_VAL;
wire [15:0] SP_VAL;

wire [15:0] INSTR_FROM_MEMORY;
wire [15:0] CURRENT_INSTR;
wire [5:0] CURRENT_INSTR_OPCODE;
wire CURRENT_INSTR_REG_ADDR;
wire [1:0] CURRENT_INSTR_REG_ADDRESS_STACK;
wire [8:0] CURRENT_INSTR_IMM;
wire [9:0] CURRENT_INSTR_BA;
wire FACT;
wire FACT_END;
wire signed [15:0] ALU_RES;
wire [3:0] ALU_FLAGS;
wire ZERO_FLAG, NEGATIVE_FLAG, CARRY_FLAG, OVERFLOW_FLAG;
wire [15:0] Extended_IMMEDIATE;
wire [15:0] Extended_BRANCH_ADDRESS;
wire [15:0] REG_INPUT;
wire [15:0] DM_INPUT;
wire [8:0] DM_ADDRESS;
wire [15:0] DM_OUT;
wire [15:0] PC_INPUT;
ProgramCounter PC(.IN(PC_INPUT),.CLK(CLK),.RST(RST), .BRA(BRA), .POP(POP), .FACT(FACT), .EN((SEL_PC & !STORE) | (BRA & ~COND_BRA) | (COND_BRA & BRZ & ZERO_FLAG) | (COND_BRA & BRN & NEGATIVE_FLAG) | (COND_BRA & BRC & CARRY_FLAG) | (COND_BRA & BRO & OVERFLOW_FLAG)),.OUT(PC_VAL));
InstructionMemory IM(.ADDRESS(PC_VAL[9:0]),.RST(RST),.OUT(INSTR_FROM_MEMORY));
InstructionRegister IR(.IN(INSTR_FROM_MEMORY),.CLK(CLK),.RST(RST),.EN(1'd1),.OUT(CURRENT_INSTR),.OPCODE(CURRENT_INSTR_OPCODE),.REGISTER_ADDRESS(CURRENT_INSTR_REG_ADDR),.REGISTER_ADDRESS_STACK(CURRENT_INSTR_REG_ADDRESS_STACK),.IMMEDIATE(CURRENT_INSTR_IMM),.BA(CURRENT_INSTR_BA));
ControlUnit CU(.OPCODE(CURRENT_INSTR_OPCODE),.REGISTER_ADDRESS(CURRENT_INSTR_REG_ADDR),.REGISTER_ADDRESS_STACK(CURRENT_INSTR_REG_ADDRESS_STACK),.IMMEDIATE(CURRENT_INSTR_IMM),.CLK(CLK),.RST(RST),.ALU(ALU),.BRA(BRA),.COND_BRA(COND_BRA),.BRZ(BRZ),.BRN(BRN),.BRC(BRC),.BRO(BRO),.LOAD(LOAD),.STORE(STORE),.COPY(COPY),.PUSH(PUSH),.POP(POP),.MOV(MOV),.SEL_FLAG(SEL_FLAG),.SEL_ACC(SEL_ACC),.SEL_X(SEL_X),.SEL_Y(SEL_Y),.SEL_PC(SEL_PC),.FACT(FACT), .FACT_END(FACT_END));
Acumulator ACC(.IN(REG_INPUT),.CLK(CLK),.RST(RST),.EN(SEL_ACC & !STORE),.OUT(ACC_VAL));
X XRegister(.IN(REG_INPUT),.CLK(CLK),.RST(RST),.EN(SEL_X & !STORE),.OUT(X_VAL));
Y YRegister(.IN(REG_INPUT),.CLK(CLK),.RST(RST),.EN(SEL_Y & !STORE),.OUT(Y_VAL));
MUX_WRITE_REG WriteDeciderRegister(.ALU_INPUT(ALU_RES),.MOV_INPUT(Extended_IMMEDIATE),.DM_INPUT(DM_OUT),.ACC_COPY(ACC_VAL),.ALU(ALU),.MOV(MOV),.LOAD(LOAD),.COPY(COPY),.IN(REG_INPUT));
ALU ArithmeticLogicUnit(.ACC(ACC_VAL),.X(X_VAL),.Y(Y_VAL),.IMMEDIATE(Extended_IMMEDIATE),.fact_reg(factorialModule.fact_OUT),.fact_val({ {7{1'b0}}, factorialModule.current_iteration[8:0] }),.OPCODE(CURRENT_INSTR_OPCODE),.EN(ALU),.CLK(CLK),.RST(RST),.REGISTER_ADDRESS(CURRENT_INSTR_REG_ADDR),.res(ALU_RES),.flags(ALU_FLAGS));
flags FlagsRegister(.IN(ALU_FLAGS),.CLK(CLK),.RST(RST),.ED(SEL_FLAG),.ZERO(ZERO_FLAG),.NEGATIVE(NEGATIVE_FLAG),.CARRY(CARRY_FLAG),.OVERFLOW(OVERFLOW_FLAG));
SignalExtender9x16 ImmediateExtender(.IN(CURRENT_INSTR_IMM),.OUT(Extended_IMMEDIATE));
REG_MUX_DM_INPUT DataMemoryInputDecider(.X(X_VAL),.Y(Y_VAL),.ACC(ACC_VAL),.PC(PC_VAL),.SEL_X(SEL_X),.SEL_Y(SEL_Y),.SEL_ACC(SEL_ACC),.SEL_PC(SEL_PC),.STORE(STORE),.IN(DM_INPUT));
DataMemory DM(.IN(DM_INPUT),.ADDR(DM_ADDRESS),.CLK(CLK),.RST(RST),.ED(STORE),.OUT(DM_OUT));
StackPointer SP(.CLK(CLK),.RST(RST),.INC(POP),.DEC(PUSH),.OUT(SP_VAL));
REG_MUX_DM_ADDR DataMemoryAddressDecider(.IMMEDIATE(CURRENT_INSTR_IMM),.SP(SP_VAL[8:0]),.LOAD(LOAD),.STORE(STORE),.PUSH(PUSH),.POP(POP),.IN(DM_ADDRESS));
BitConverter10x16 BranchAddressExtender(.IN(CURRENT_INSTR_BA),.OUT(Extended_BRANCH_ADDRESS));
ProgramCounterInputDecider PCInputDecider(.POPInput(REG_INPUT),.BRAInput(Extended_BRANCH_ADDRESS),.POP(POP),.BRA(BRA),.ProgramCounterInput(PC_INPUT)); 

endmodule